-- Universidade Federal de Minas Gerais
-- Escola de Engenharia
-- Departamento de Engenharia Eletrônica
-- Autoria: Professor Ricardo de Oliveira Duarte
-- Unidade de controle ciclo único (look-up table) do processador
-- puramente combinacional
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- unidade de controle
entity unidade_de_controle_ciclo_unico is
    generic (
        INSTR_WIDTH       : natural := 16;
        OPCODE_WIDTH      : natural := 5;
        DP_CTRL_BUS_WIDTH : natural := 17;
        ULA_CTRL_WIDTH    : natural := 3
    );
    port (
        instrucao : in std_logic_vector(INSTR_WIDTH - 1 downto 0);       -- instrução
        controle  : out std_logic_vector(DP_CTRL_BUS_WIDTH - 1 downto 0); -- controle da via
        in_flag_zero : in std_logic
    );
end unidade_de_controle_ciclo_unico;

architecture beh of unidade_de_controle_ciclo_unico is
    -- As linhas abaixo não produzem erro de compilação no Quartus II, mas no Modelsim (GHDL) produzem.	
    --signal inst_aux : std_logic_vector (INSTR_WIDTH-1 downto 0);			-- instrucao
    --signal opcode   : std_logic_vector (OPCODE_WIDTH-1 downto 0);			-- opcode
    --signal ctrl_aux : std_logic_vector (DP_CTRL_BUS_WIDTH-1 downto 0);		-- controle

    signal inst_aux : std_logic_vector (15 downto 0); -- instrucao
    signal opcode   : std_logic_vector (4 downto 0);  -- opcode
    signal ctrl_aux : std_logic_vector (16 downto 0);  -- controle

begin
    inst_aux <= instrucao;
    -- A linha abaixo não produz erro de compilação no Quartus II, mas no Modelsim (GHDL) produz.	
    --	opcode <= inst_aux (INSTR_WIDTH-1 downto INSTR_WIDTH-OPCODE_WIDTH);
    opcode <= inst_aux (4 downto 0);

    -- UL UL UL MA1 MD1 MLM WE1 WE2 RA RB MA MB WEData RDData MPC MPC PCW
    -- 0  1  2  3   4   5   6   7   8  9  10 11 12     13     14  15  16

    process (opcode)
    begin
        case opcode is
                -- NAND	
            when "00000" =>
                ctrl_aux <= "00000000000000000";
                -- OR
            when "00001" =>
                ctrl_aux <= "00000000000000000";
                -- ADD
            when "00010" =>
                ctrl_aux <= "00000000000000000";
                -- SUB	
            when "00100" =>
                ctrl_aux <= "00000000000000000";
                -- XOR
            when "01100" =>
                ctrl_aux <= "00000000000000000";
            when others =>
                ctrl_aux <= (others => '0');
        end case;
    end process;
    controle <= ctrl_aux;
end beh;